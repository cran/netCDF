netcdf panom {
dimensions:
	XPCIPSEAS1_73 = 73 ;
	YPCIPSEAS1_37 = 37 ;
variables:
	double XPCIPSEAS1_73(XPCIPSEAS1_73) ;
		XPCIPSEAS1_73:units = "degrees_east" ;
		XPCIPSEAS1_73:modulo = " " ;
		XPCIPSEAS1_73:point_spacing = "even" ;
	double YPCIPSEAS1_37(YPCIPSEAS1_37) ;
		YPCIPSEAS1_37:units = "degrees_north" ;
		YPCIPSEAS1_37:point_spacing = "even" ;
	float PANOM(YPCIPSEAS1_37, XPCIPSEAS1_73) ;
		PANOM:missing_value = -9999.99f ;
		PANOM:_FillValue = -9999.99f ;
		PANOM:long_name = "Seasonal precip anomaly" ;
		PANOM:long_name_mod = "T=15-JAN-1989@ITP" ;
		PANOM:history = "From land_precip" ;
		PANOM:units = "mm" ;

// global attributes:
		:history = "FERRET V4.91 (PMEL v4.91b3/GUI) 27-Dec-99" ;
data:

 XPCIPSEAS1_73 = 0, 5, 10, 15, 20, 25, 30, 35, 40, 45, 50, 55, 60, 65, 70, 
    75, 80, 85, 90, 95, 100, 105, 110, 115, 120, 125, 130, 135, 140, 145, 
    150, 155, 160, 165, 170, 175, 180, 185, 190, 195, 200, 205, 210, 215, 
    220, 225, 230, 235, 240, 245, 250, 255, 260, 265, 270, 275, 280, 285, 
    290, 295, 300, 305, 310, 315, 320, 325, 330, 335, 340, 345, 350, 355, 360 ;

 YPCIPSEAS1_37 = -62, -58, -54, -50, -46, -42, -38, -34, -30, -26, -22, -18, 
    -14, -10, -6, -2, 2, 6, 10, 14, 18, 22, 26, 30, 34, 38, 42, 46, 50, 54, 
    58, 62, 66, 70, 74, 78, 82 ;

 PANOM =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, -60.83994, _, 83.0585, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 37.76834, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 9.44264, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, -250.91, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 6.415421, _, _, -66.5342, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -17.49778, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, -23.92323, -20.62855, _, _, _, -108.904, 63.99384, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -46.99278, 
    -19.25145, -34.19439, _, _, _, _, _, _, _, _, _, _, -110.0103, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, -20.16297, 9.24453, 63.13947, _, _, _, _, 123.3779, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -132.0978, -29.74171, 
    -70.87589, -55.7188, -10.76826, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, -13.08612, -47.37563, -89.76459, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 69.19541, -3.252753, _, _, -3.57578, -23.05547, 
    7.318983, 28.0409, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, -43.12314, _, 15.42809, -127.507, -4.317777, 
    -45.79231, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 17.61214, 53.78723, 78.82139, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 26.81602, 27.16825, 73.86526, 65.20012, 7.829914, 
    15.56462, -48.72092, -60.39011, 121.7619, 16.44221, _, 8.585036, _, 
    230.3234, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    -0.9855256, -79.28306, -122.7436, -125.6138, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, 29.01458, -65.77568, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, -21.22568, 32.91608, _, _, _, -29.81698, -132.3066, -18.80531, 
    169.4789, _, _, _, _, _, _, _, _, _, _, _, -74.25889, _, _, _, _, _, _, 
    -112.7924, _, _, _, _, _, _, _, _, -368.6052, -60.58345, -9.9859, 
    128.4334, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, -91.82261, -136.3947, _, 38.89001, _, _, 15.68039, _, _, 
    _, _, _, _, _, _, _, _, -65.89575, 78.64118, _, _, -56.2993, _, 
    -57.16877, 15.16337, _, _, 293.3743, _, _, _, _, _, _, _, _, -124.2698, 
    _, _, -160.5811, _, _, _, _, _, _, _, _, _, _, _, _, -0.05098506, 
    65.79301, -73.38407, _, _, -112.7564, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, 118.8562, 58.21017, 60.72109, _, 193.4481, -58.49446, _, 
    50.16521, -98.53196, _, _, _, _, _, _, _, _, _, _, -196.5944, -172.3974, 
    -177.8775, _, -187.2111, -260.6529, -173.2925, _, _, _, _, _, 697.7068, 
    _, _, _, _, _, -207.8741, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    0.8373526, _, 27.37533, _, _, _, _, _, _, _, _, _, _, -77.7636, _,
  _, _, _, _, _, _, 7.259945, 171.4049, -21.69259, 377.8698, 310.3261, _, _, 
    _, _, _, _, _, _, 44.11475, _, _, _, _, _, _, -137.2703, -101.001, 
    86.95312, -0.4078361, _, _, _, _, _, _, _, 216.3532, 379.7586, _, _, _, 
    _, -177.0526, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    193.2924, _, -79.22112, 79.3955, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, -85.06818, _, _, _, _, 294.688, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 117.4031, 276.1908, _, _, _, _, _, _, _, -226.1997, 
    _, _, _, _, _, _, _, -34.44004, _, _, _, _, _, _, _, _, _, _, _, _, 
    -143.2069, _, _, _, _, -96.3312, _, -16.57234, 29.85958, _, _, _, _, _, 
    _, _,
  _, _, _, 110.5388, _, _, _, 40.4399, 175.8595, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, -2.0407, _, _, _, _, _, _, _, 
    -85.29628, _, _, _, _, _, _, _, _,
  _, _, _, -143.881, _, _, 156.8751, 50.36941, 47.65427, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, -157.8435, _, _, 204.3818, _, 
    _, 445.2486, _, 250.9173, _, 82.70246, _, _, _, _, _, _, _, _,
  _, _, -88.12541, -134.525, _, _, _, _, 38.47545, _, _, _, _, _, _, _, _, _, 
    _, _, -50.14315, -390.7137, 150.5068, 202.3315, _, _, _, _, _, _, _, _, 
    _, _, _, -659.4767, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  -8.640877, _, -63.45637, 10.12378, -35.59931, _, _, _, _, _, _, _, _, _, _, 
    _, -165.8574, _, _, _, -151.3594, _, _, 9.801895, -95.5917, _, _, 
    356.9156, _, _, -65.14896, _, 183.2258, _, 83.17491, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -24.27607, 3.587367, _, 
    277.3524, 872.5285, _, _, _, _, _, _, _, -80.79266, -70.43465, -8.640877,
  -8.827262, -3.237782, _, 3.67062, -1.257576, _, _, _, -21.99358, 14.70745, 
    _, _, _, _, _, -10.1776, -155.9246, _, _, -102.7759, -125.4791, _, _, _, 
    _, 248.279, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, -2.392779, -5.816735, 62.41625, _, _, 
    _, _, _, _, _, _, -47.73812, -50.58704, -6.212092, -8.827262,
  -1.341473, -0.1906632, -0.2911037, -0.009983227, -0.1911141, -0.01820234, 
    0.01382935, -0.01252876, _, _, _, _, _, _, _, -3.696085, -60.63747, _, _, 
    _, -9.879082, -42.91717, _, _, -29.16268, 458.3217, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 192.5159, 
    15.5261, _, _, 106.5822, _, _, _, _, _, _, _, _, _, _, -1.735779, 
    -1.513345, -0.9069598, -1.341473,
  _, _, -0.1486886, -0.3126243, _, _, -0.1794998, -0.07272431, _, _, _, 
    -7.399639, _, _, _, 1.333859, -8.477449, -40.84721, _, _, -26.23489, 
    -29.50096, _, _, -23.81884, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 317.1124, _, _, _, _, _, _, _, _, _, _, _, -11.01943, 24.16735, _, _, 
    156.618, 200.218, 46.16806, _, _, _, _, _, _, _, _, _, -3.217111, 
    -2.927739, -0.6604142, _,
  _, -5.170388, _, _, _, _, _, _, _, _, _, _, -14.97013, _, 2.336949, 
    -17.23391, -39.93641, _, -22.23516, _, _, _, -4.107807, 39.24355, 
    -319.1222, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 226.6151, _, _, 
    _, _, _, _, _, _, _, _, -7.56452, _, _, 229.392, _, 88.74849, _, _, _, _, 
    _, _, _, _, _, _, _, _, -9.800809, _, _, _,
  _, _, -6.648261, _, _, _, _, _, _, -32.95912, -42.93214, _, _, -41.49984, 
    -8.141667, -5.430104, _, 11.11928, 21.11701, 43.54676, -53.59657, 
    -35.10037, -9.56853, _, _, -267.7061, -167.3801, _, -29.85413, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -11.22547, 
    -77.2644, -49.1427, _, _, -87.02564, -57.67956, _, _, _, _, _, _, _, _, 
    _, _, _, _, -4.231858, -8.700909, _,
  _, _, _, -26.36925, _, _, _, -12.57852, _, _, _, _, _, -21.64325, 
    -16.49421, 18.67676, _, _, -3.314471, -3.997028, _, 7.069686, _, 91.9242, 
    13.7243, _, -108.106, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, -54.38895, -32.63589, 9.835123, 73.12362, -99.47884, 
    -172.3376, -162.073, -89.62088, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    -78.28036, 63.46296, _,
  _, -26.72347, 8.805434, -44.56263, _, -158.3662, -35.20942, -6.674884, _, 
    _, _, _, _, _, -33.03755, 47.47972, _, _, _, _, _, _, 44.51365, 59.78323, 
    _, 1172.558, 129.3317, 161.8324, -19.16572, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, -95.39229, -5.306077, -36.23935, -4.965796, 
    12.83724, 7.305501, 204.35, -116.99, -122.9376, -153.2392, _, _, _, _, _, 
    _, _, _, _, _, _, _, -93.80145, -67.12103, _,
  -1.717584, -118.7088, -56.38537, _, -412.8006, -54.31877, -141.7158, 
    -76.71363, -100.5024, -0.8512377, _, _, -20.98711, _, _, -9.547184, _, _, 
    _, _, -2.093194, 12.40598, _, 7.388703, _, 30.3397, 263.2059, -133.0448, 
    -47.89138, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    -333.3784, -56.67388, -13.51546, -3.462934, 15.79743, -25.7073, 
    -2.266124, 53.98174, 145.1199, -85.73612, -88.96214, _, _, _, _, _, _, _, 
    _, -169.4139, -12.80225, _, _, -113.493, -118.9219, -1.717584,
  -10.36692, -96.99019, -94.21998, -193.0862, -297.1182, -134.376, -48.50313, 
    -13.17763, -176.3069, -42.06554, _, 2.139189, 21.28618, _, -8.247773, 
    40.4493, _, _, 5.066395, -4.235467, _, -3.680508, _, _, _, -7.565632, 
    -5.060678, _, -48.69943, -84.15612, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, -354.6175, -53.79551, -40.50053, -10.70428, -7.937628, 
    -3.614027, -8.183489, -38.49168, -30.78896, -41.02889, -79.147, 
    -160.2718, -124.1284, _, _, _, _, _, _, _, _, _, _, -179.139, -53.63588, 
    -10.36692,
  -85.34901, -14.31164, -36.65707, -104.2277, -52.93326, -25.64645, 
    -14.94428, -0.3847288, 25.36914, 17.87424, 12.38775, _, _, _, _, 
    27.66035, -9.546387, _, _, -1.809758, _, -0.1253024, 1.210593, _, _, _, 
    _, _, -109.8757, -47.16254, -63.73768, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, -254.9716, -21.26587, -35.75864, 22.50956, -1.594979, 
    5.582354, -2.908544, 0.4468629, 14.9008, 13.99885, -69.71013, -83.835, 
    -73.15734, -65.6779, -43.536, _, _, _, _, _, _, _, _, _, -44.70679, 
    -85.34901,
  _, -25.05503, 0.909149, 4.068902, -15.48613, -15.55287, 10.73156, 
    -23.00594, 11.09395, -8.73, _, 8.66159, _, 41.12492, _, 29.62023, 
    4.350735, _, _, _, -0.3921933, -1.735978, _, _, 51.6199, _, -3.855187, 
    52.25793, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    -181.2617, -77.27795, -4.327448, 31.73302, 4.876374, 7.603703, -14.7129, 
    8.450061, 11.65311, _, -3.642859, _, -34.66219, -54.93539, -77.7609, 
    38.2627, _, _, _, _, _, _, _, _, -26.13617, -62.86872, _,
  _, -44.13643, -32.09285, -39.18492, -9.496386, 2.467873, 17.80319, _, 
    55.40229, _, 54.07602, _, _, 17.40899, _, 50.69022, _, 5.16944, 
    -5.470432, _, _, 1.38095, _, -2.158989, _, _, 70.44788, _, 0.2454958, _, 
    _, _, 179.6815, _, _, -27.38231, _, _, _, 94.39591, _, _, _, _, _, 
    37.31007, -115.8227, -2.901906, -27.33115, -19.72387, -11.60584, 
    -27.04964, -15.44787, _, 0.008716182, _, _, _, _, _, -137.0221, _, _, _, 
    _, _, _, _, _, _, 54.21545, -34.36502, _,
  _, 159.7191, -25.29827, -4.511099, -42.35978, _, 16.15592, _, 3.932329, _, 
    45.46205, _, 21.97366, _, 19.75354, _, _, 19.7237, 6.232504, -5.935946, 
    -17.6826, _, 4.21204, _, _, 54.73153, _, _, _, 19.3385, _, _, _, _, _, _, 
    _, _, 81.65874, _, _, 3.369525, -24.1306, _, 203.8421, -24.85327, 
    36.90949, -25.72957, -28.04343, _, -18.45171, _, _, 7.735264, _, _, 
    10.76833, _, -44.67204, _, _, _, _, _, _, _, _, _, _, _, _, 186.3948, _,
  _, _, 88.7947, -4.68189, 0.3717763, 62.6705, 76.30644, _, _, _, _, _, _, _, 
    25.50847, _, _, _, 44.56701, _, _, _, -8.477483, _, 45.34235, _, 
    19.24039, _, _, 3.095733, -20.59076, _, _, 53.12723, _, _, _, _, _, _, 
    52.68505, 73.62836, 2.171958, 12.9189, -10.13364, -16.1688, -28.22514, _, 
    _, -11.51267, -26.43181, _, _, _, _, _, _, _, -39.68225, _, _, _, _, _, 
    _, _, _, _, _, _, _, 296.1394, _,
  _, _, _, 145.04, _, 40.51064, 55.22863, _, 49.25991, _, _, _, _, 18.84679, 
    _, _, _, _, 33.09284, _, 11.29396, _, _, _, _, _, _, 18.53217, _, _, 
    -11.94572, _, _, _, 21.73841, _, 144.2157, _, 8.242409, 43.477, _, _, 
    38.7971, 21.64352, _, _, _, -0.6746025, _, 6.676734, _, _, _, 9.826651, 
    _, -20.56243, _, _, _, _, _, _, -24.07618, _, -46.29916, _, _, 141.1345, 
    169.1395, -29.23124, _, _, _,
  _, _, _, _, 171.9912, 45.65324, 159.3972, 11.77927, _, 5.567222, _, _, _, 
    _, _, -20.83051, _, _, _, _, _, _, 1.146449, _, _, _, _, _, _, _, 
    -2.567884, _, -13.05538, _, _, _, -6.481011, _, _, _, _, 0.9754165, _, _, 
    _, _, _, _, _, _, _, 4.443224, _, _, _, _, _, _, -8.773625, _, _, 
    -18.63514, _, _, _, _, _, _, -68.78065, _, 86.3035, _, _,
  _, _, _, _, 55.16798, _, _, _, _, _, _, _, _, _, _, _, 39.34165, _, _, _, 
    _, 1.186213, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, -3.593647, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -20.23678, _, _, _, _, _, 
    -13.4397, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 16.92883, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, -13.8899, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 9.575752, _, _, _, _, 15.66923, _, _, _, _, _, _, _, _, 
    _, _, _, _ ;
}
