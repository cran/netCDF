netcdf x {
dimensions:
        x = 3 ;
        y = 4 ;
variables:
        float x(x, y) ;
data:

 x =
  1, 2, 3, 4,
  5, 6, 7, 8,
  9, 10, 11, 12 ;
}
